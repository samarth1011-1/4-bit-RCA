module rca()
endmodule